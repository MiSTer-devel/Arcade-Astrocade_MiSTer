library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity BALLY_STARPOS is
  port (
    ADDR        : in    std_logic_vector(9 downto 0);
    DATA        : out   std_logic_vector(8 downto 0)
    );
end;

-- Horizontal star positions, X"160" is end of that vertical trace.

-- some at bottom are probably off-screen, may tidy up later!

architecture RTL of BALLY_STARPOS is

  type ROM_ARRAY is array(0 to 563) of std_logic_vector(11 downto 0);
  constant ROM : ROM_ARRAY := (
		X"160",
		X"026",X"0BC",X"160",
		X"027",X"082",X"160",
		X"005",X"160",
		X"009",X"0AE",X"0B6",X"160",
		X"160",
		X"012",X"160",
		X"0C8",X"160",
		X"007",X"013",X"160",
		X"0E1",X"102",X"160",
		X"160",
		X"072",X"160",
		X"160",
		X"0EE",X"160",
		X"08C",X"160",
		X"0D7",X"160",
		X"038",X"0A5",X"160",
		X"160",
		X"114",X"160",
		X"160",
		X"0A8",X"160",
		X"0D0",X"160",
		X"160",
		X"160",
		X"055",X"05D",X"11B",X"160",
		X"026",X"051",X"160",
		X"02E",X"0FA",X"139",X"160",
		X"12F",X"160",
		X"072",X"11C",X"160",
		X"12D",X"160",
		X"004",X"036",X"160",
		X"021",X"0C4",X"160",
		X"160",
		X"160",
		X"09F",X"12B",X"160",
		X"12F",X"160",
		X"160",
		X"0FC",X"160",
		X"160",
		X"160",
		X"160",
		X"160",
		X"066",X"160",
		X"023",X"160",
		X"020",X"160",
		X"07B",X"087",X"160",
		X"00A",X"01F",X"0AD",X"160",
		X"135",X"160",
		X"0C0",X"160",
		X"114",X"160",
		X"0EE",X"160",
		X"0F9",X"160",
		X"0B7",X"160",
		X"02F",X"0AC",X"160",
		X"021",X"160",
		X"118",X"160",
		X"0A0",X"0D1",X"0E5",X"160",
		X"098",X"122",X"160",
		X"113",X"160",
		X"031",X"0F6",X"160",
		X"160",
		X"06B",X"160",
		X"160",
		X"0A9",X"160",
		X"051",X"160",
		X"0EB",X"160",
		X"0C3",X"160",
		X"11B",X"160",
		X"095",X"0DC",X"160",
		X"160",
		X"160",
		X"0AF",X"102",X"13F",X"160",
		X"04B",X"0BB",X"10B",X"160",
		X"0C8",X"160",
		X"0DF",X"160",
		X"027",X"033",X"160",
		X"006",X"160",
		X"0B8",X"0F2",X"12A",X"160",
		X"138",X"160",
		X"160",
		X"01F",X"160",
		X"069",X"160",
		X"160",
		X"058",X"10F",X"160",
		X"160",
		X"040",X"09F",X"160",
		X"0E4",X"112",X"160",
		X"160",
		X"044",X"160",
		X"00D",X"0E4",X"160",
		X"01C",X"0CE",X"120",X"160",
		X"134",X"160",
		X"00A",X"079",X"134",X"160",
		X"08F",X"0E4",X"160",
		X"124",X"160",
		X"008",X"0A4",X"160",
		X"003",X"133",X"160",
		X"109",X"160",
		X"022",X"041",X"0B2",X"0E4",X"0F8",X"112",X"128",X"134",X"160",
		X"0CC",X"116",X"160",
		X"03B",X"160",
		X"160",
		X"10E",X"160",
		X"04A",X"160",
		X"0CD",X"160",
		X"135",X"160",
		X"160",
		X"0F1",X"160",
		X"007",X"060",X"160",
		X"124",X"160",
		X"11B",X"160",
		X"160",
		X"06D",X"0E7",X"12A",X"160",
		X"00B",X"09B",X"111",X"160",
		X"160",
		X"024",X"0E0",X"160",
		X"160",
		X"016",X"093",X"160",
		X"160",
		X"027",X"0CE",X"0FF",X"160",
		X"0CC",X"160",
		X"160",
		X"0FA",X"160",
		X"09A",X"0A6",X"160",
		X"03E",X"160",
		X"085",X"160",
		X"089",X"116",X"160",
		X"033",X"09B",X"160",
		X"160",
		X"017",X"109",X"160",
		X"043",X"160",
		X"0CB",X"102",X"160",
		X"07C",X"160",
		X"0AA",X"160",
		X"0AE",X"160",
		X"096",X"160",
		X"07B",X"12B",X"160",
		X"0AF",X"160",
		X"13B",X"160",
		X"00E",X"160",
		X"160",
		X"160",
		X"053",X"160",
		X"160",
		X"006",X"0B5",X"0FC",X"160",
		X"160",
		X"072",X"0B4",X"160",
		X"03F",X"160",
		X"018",X"160",
		X"06D",X"160",
		X"044",X"078",X"0D6",X"12F",X"160",
		X"036",X"0FB",X"114",X"160",
		X"02B",X"160",
		X"160",
		X"0B5",X"160",
		X"01F",X"0EF",X"11B",X"160",
		X"0A1",X"104",X"160",
		X"076",X"160",
		X"048",X"075",X"0DD",X"160",
		X"160",
		X"0CE",X"160",
		X"0F0",X"160",
		X"009",X"028",X"160",
		X"160",
		X"022",X"056",X"160",
		X"042",X"0D2",X"160",
		X"0F5",X"160",
		X"05B",X"160",
		X"13F",X"160",
		X"0A7",X"160",
		X"081",X"134",X"160",
		X"0D8",X"160",
		X"047",X"160",
		X"015",X"05E",X"160",
		X"05D",X"160",
		X"160",
		X"037",X"160",
		X"0B7",X"119",X"160",
		X"160",
		X"0DA",X"160",
		X"032",X"10A",X"160",
		X"028",X"160",
		X"08E",X"160",
		X"0B5",X"160",
		X"0B3",X"160",
		X"00A",X"129",X"160",
		X"124",X"160",
		X"028",X"160",
		X"063",X"160",
		X"076",X"160",
		X"160",
		X"082",X"0C7",X"0F4",X"160",
		X"160",
		X"068",X"160",
		X"02A",X"160",
		X"0B2",X"0E9",X"160",
		X"160",
		X"031",X"077",X"091",X"0A7",X"0B3",X"160",
		X"04B",X"095",X"0EB",X"160",
		X"160",
		X"160",
		X"08D",X"10D",X"160",
		X"06E",X"160",
		X"04C",X"160",
		X"0B4",X"0FC",X"160",
		X"01E",X"0CC",X"0D8",X"160",
		X"070",X"160",
		X"160",
		X"079",X"0A3",X"0E3",X"160",
		X"09A",X"160",
		X"028",X"09B",X"160",
		X"026",X"066",X"160",
		X"090",X"09C",X"160",
		X"034",X"0B5",X"0FD",X"160",
		X"05F",X"0C6",X"160",
		X"0CE",X"160",
		X"012",X"08D",X"160",
		X"0AD",X"112",X"160",
		X"160",
		X"160",
		X"160",
		X"160",
		X"160",
		X"160",
		X"160",
		X"160",
		X"160",
		X"160",
		X"160",
		X"160",
		X"160",
		X"160",
		X"160",
		X"160",
		X"160",
		X"160",
		X"160",
		X"160",
		X"160",
		X"160",
		X"160",
		X"100",X"160",
		X"0CF",X"160",
		X"034",X"04D",X"160",
		X"160",
		X"160",
		X"075",X"160",
		X"160",
		X"135",X"160",
		X"0AE",X"160",
		X"160",
		X"160",
		X"04A",X"160",
		X"0F1",X"160",
		X"06E",X"160",
		X"020",X"083",X"160",
		X"160",
		X"0B8",X"135",X"160",
		X"160",
		X"04D",X"160",
		X"160",
		X"018",X"08E",X"0EB",X"160",
		X"160",
		X"FFF" -- End Marker
);

begin

  p_rom : process(ADDR)
  begin
     DATA <= ROM(to_integer(unsigned(ADDR)))(8 downto 0);
  end process;

end RTL;

